`timescale 1ns / 1ps
//Image generation part
module Video_Generator(
    input clk,
    input [11:0]bpos_x,
    input [11:0]bpos_y,
    input [11:0]pippos0_x1,
    input [11:0]pippos0_y1,
    input [11:0]pippos0_x2,
    input [11:0]pippos0_y2,
    input [11:0]pippos1_x1,
    input [11:0]pippos1_y1,
    input [11:0]pippos1_x2,
    input [11:0]pippos1_y2,
    input [11:0]pippos2_x1,
    input [11:0]pippos2_y1,
    input [11:0]pippos2_x2,
    input [11:0]pippos2_y2,
    input start_num0,
    input start_num1,
    input start_num2,
	input [4:0]point1,
	input [4:0]point2,
	input [4:0]point3,
	input game_over,
    input RGB_VDE,
    input [11:0]Set_X,
    input [11:0]Set_Y,
    output reg[23:0]RGB_Data=24'hffff00    //RBG
    );
    reg [11:0]Address=0;
    reg [255:0] rom_data0 = 256'h00000000000007E01818381C300C300C300C300C300C38181C1007E000000000;
    reg [255:0] rom_data1 = 256'h00000000000000800780018001800180018001800180018001800FF800000000;
    reg [255:0] rom_data2 = 256'h0000000000000FF03018380C101800180060018006000804300C3FF800000000;
    reg [255:0] rom_data3 = 256'h0000000000000FE0301838180018006001F00018000C380C30180FE000000000;
    reg [255:0] rom_data4 = 256'h000000000000003000F0017002700C70107020707FFE0070007003FE00000000;
    reg [255:0] rom_data5 = 256'h0000000000001FF810001000100017F01818000C000C380C30180FE000000000;
    reg [255:0] rom_data6 = 256'h00000000000007F008181000300037F0380C300C300C300C181807E000000000;
    reg [255:0] rom_data7 = 256'h0000000000001FFC300820100020004000800180030003000380030000000000;
    reg [255:0] rom_data8 = 256'h0000000000000FF03008300C38080F300DE03038600C600C30080FF000000000;
    reg [255:0] rom_data9 = 256'h0000000000000FE03018300C700C301C382C0FCC001C001838300FC000000000;
    
    reg [15:0] char_0_r [15:0] ;
    reg [15:0] char_1_r [15:0] ;
    reg [15:0] char_2_r [15:0] ;
    reg [15:0] char_3_r [15:0] ;
    reg [15:0] char_4_r [15:0] ;
    reg [15:0] char_5_r [15:0] ;
    reg [15:0] char_6_r [15:0] ;
    reg [15:0] char_7_r [15:0] ;
    reg [15:0] char_8_r [15:0] ;
    reg [15:0] char_9_r [15:0] ;
    
    wire [23:0]bird_data;
	//wire Num_Data;
    // wire [7:0]R_Data;
    // wire [7:0]G_Data;
    // wire [7:0]B_Data;

always@(*)
        begin
           
			// if(Set_X>=12'd720&&Set_X<=12'd780&&Set_Y>=12'd360&&Set_Y<=12'd400)
			//  begin  Address<=(Set_Y-12'd359)*40+(Set_X-12'd719);RGB_Data<={bird_data[23:16],bird_data[7:0],bird_data[15:8]};  end
            if(Set_X<=12'd1280&&Set_X>=12'd0&&Set_Y<=12'd720&&Set_Y>=12'd0&&game_over)
			   begin RGB_Data<=24'hed869b; end
			else if ( (Set_X>=bpos_x-12'd30) && (Set_X<=bpos_x+12'd30) &&(Set_Y>=bpos_y-12'd20)&&(Set_Y<=bpos_y+12'd20))
               begin
                  RGB_Data<=24'h86edb0;
               end
			// else if ( (Set_X>=12'd1100) && (Set_X<=12'd1140) &&(Set_Y>=12'd0)&&(Set_Y<=12'd40))
            //    begin
            //       if(game_over) RGB_Data<=24'hed869b;
			// 	  else RGB_Data<=24'h7558ff;
            //    end
            else if(Set_X>=12'd1000&&Set_X<=12'd1015&&Set_Y>=12'd0&&Set_Y<=12'd15)
                begin
                   case(point1)
				     4'd0: RGB_Data<=char_0_r[Set_Y][12'd984-Set_X]?24'h20ffb2:24'hffbffa;
				     4'd1: RGB_Data<=char_1_r[Set_Y][12'd984-Set_X]?24'h20ffb2:24'hffbffa;
				     4'd2: RGB_Data<=char_2_r[Set_Y][12'd984-Set_X]?24'h20ffb2:24'hffbffa;
				     4'd3: RGB_Data<=char_3_r[Set_Y][12'd984-Set_X]?24'h20ffb2:24'hffbffa;
				     4'd4: RGB_Data<=char_4_r[Set_Y][12'd984-Set_X]?24'h20ffb2:24'hffbffa;
				     4'd5: RGB_Data<=char_5_r[Set_Y][12'd984-Set_X]?24'h20ffb2:24'hffbffa;
				     4'd6: RGB_Data<=char_6_r[Set_Y][12'd984-Set_X]?24'h20ffb2:24'hffbffa;
				     4'd7: RGB_Data<=char_7_r[Set_Y][12'd984-Set_X]?24'h20ffb2:24'hffbffa;
				     4'd8: RGB_Data<=char_8_r[Set_Y][12'd984-Set_X]?24'h20ffb2:24'hffbffa;
				     4'd9: RGB_Data<=char_9_r[Set_Y][12'd984-Set_X]?24'h20ffb2:24'hffbffa;
				     default: RGB_Data<=char_0_r[Set_Y][12'd984-Set_X]?24'h20ffb2:24'hffbffa;
				   endcase
                end
			else if(Set_X>=12'd984&&Set_X<=12'd999&&Set_Y>=12'd0&&Set_Y<=12'd15)
                begin
                   case(point2)
				     4'd0: RGB_Data<=char_0_r[Set_Y][12'd968-Set_X]?24'h20ffb2:24'hffbffa;
				     4'd1: RGB_Data<=char_1_r[Set_Y][12'd968-Set_X]?24'h20ffb2:24'hffbffa;
				     4'd2: RGB_Data<=char_2_r[Set_Y][12'd968-Set_X]?24'h20ffb2:24'hffbffa;
				     4'd3: RGB_Data<=char_3_r[Set_Y][12'd968-Set_X]?24'h20ffb2:24'hffbffa;
				     4'd4: RGB_Data<=char_4_r[Set_Y][12'd968-Set_X]?24'h20ffb2:24'hffbffa;
				     4'd5: RGB_Data<=char_5_r[Set_Y][12'd968-Set_X]?24'h20ffb2:24'hffbffa;
				     4'd6: RGB_Data<=char_6_r[Set_Y][12'd968-Set_X]?24'h20ffb2:24'hffbffa;
				     4'd7: RGB_Data<=char_7_r[Set_Y][12'd968-Set_X]?24'h20ffb2:24'hffbffa;
				     4'd8: RGB_Data<=char_8_r[Set_Y][12'd968-Set_X]?24'h20ffb2:24'hffbffa;
				     4'd9: RGB_Data<=char_9_r[Set_Y][12'd968-Set_X]?24'h20ffb2:24'hffbffa;
				     default: RGB_Data<=char_0_r[Set_Y][12'd968-Set_X]?24'h20ffb2:24'hffbffa;
				   endcase
                end
			else if(Set_X>=12'd968&&Set_X<=12'd983&&Set_Y>=12'd0&&Set_Y<=12'd15)
			    begin
				  case(point3)
					4'd0: RGB_Data<=char_0_r[Set_Y][12'd952-Set_X]?24'h20ffb2:24'hffbffa;
					4'd1: RGB_Data<=char_1_r[Set_Y][12'd952-Set_X]?24'h20ffb2:24'hffbffa;
					4'd2: RGB_Data<=char_2_r[Set_Y][12'd952-Set_X]?24'h20ffb2:24'hffbffa;
					4'd3: RGB_Data<=char_3_r[Set_Y][12'd952-Set_X]?24'h20ffb2:24'hffbffa;
					4'd4: RGB_Data<=char_4_r[Set_Y][12'd952-Set_X]?24'h20ffb2:24'hffbffa;
					4'd5: RGB_Data<=char_5_r[Set_Y][12'd952-Set_X]?24'h20ffb2:24'hffbffa;
					4'd6: RGB_Data<=char_6_r[Set_Y][12'd952-Set_X]?24'h20ffb2:24'hffbffa;
					4'd7: RGB_Data<=char_7_r[Set_Y][12'd952-Set_X]?24'h20ffb2:24'hffbffa;
					4'd8: RGB_Data<=char_8_r[Set_Y][12'd952-Set_X]?24'h20ffb2:24'hffbffa;
					4'd9: RGB_Data<=char_9_r[Set_Y][12'd952-Set_X]?24'h20ffb2:24'hffbffa;
					default: RGB_Data<=char_0_r[Set_Y][12'd952-Set_X]?24'h20ffb2:24'hffbffa;
				endcase
			     end
            else if(( (Set_X >= pippos0_x1-12'd25 && Set_X <=pippos0_x1+12'd25 && ((Set_Y>=0 && Set_Y<=pippos0_y1)||( Set_Y>=pippos0_y2 && Set_Y<=12'd720)))
                     ||((Set_X>=pippos0_x1-12'd40&&Set_X <=pippos0_x1+12'd40)&&((Set_Y>=pippos0_y1-12'd10&&Set_Y<=pippos0_y1+12'd10)||(Set_Y>=pippos0_y2-12'd10&&Set_Y<=pippos0_y2+12'd10)))
                     )&&(start_num0))
               begin  
                   RGB_Data<= 24'h86c3ed;
               end
            else if(( (Set_X >= pippos1_x1-12'd25 && Set_X <=pippos1_x1+12'd25 && ((Set_Y>=0 && Set_Y<=pippos1_y1)||( Set_Y>=pippos1_y2 && Set_Y<=12'd720)))
                     ||((Set_X>=pippos1_x1-12'd40&&Set_X <=pippos1_x1+12'd40)&&((Set_Y>=pippos1_y1-12'd10&&Set_Y<=pippos1_y1+12'd10)||(Set_Y>=pippos1_y2-12'd10&&Set_Y<=pippos1_y2+12'd10)))
                     )&&(start_num1)) 
               begin  
                   RGB_Data<= 24'h9cd3fa;
               end
            else if(( (Set_X >= pippos2_x1-12'd25 && Set_X <=pippos2_x1+12'd25 && ((Set_Y>=0 && Set_Y<=pippos2_y1)||( Set_Y>=pippos2_y2 && Set_Y<=12'd720)))
                     ||((Set_X>=pippos2_x1-12'd40&&Set_X <=pippos2_x1+12'd40)&&((Set_Y>=pippos2_y1-12'd10&&Set_Y<=pippos2_y1+12'd10)||(Set_Y>=pippos2_y2-12'd10&&Set_Y<=pippos2_y2+12'd10)))
                     ) &&(start_num2))
               begin  
                   RGB_Data<=24'hbc9cfa;
               end   
            else
               RGB_Data<=24'hffbffa; 
         end

   bird_ROM bird_ROM0(
     .clka(clk),    // input wire clka
     .ena(1),      // input wire ena
     .addra(Address),  // input wire [13 : 0] addra
     .douta(bird_data)  // output wire [23 : 0] douta
   );
always@(posedge clk)
		begin
			char_0_r[0 ] <= rom_data0[255:240]	;
			char_0_r[1 ] <= rom_data0[239:224]	;
			char_0_r[2 ] <= rom_data0[223:208]	;
			char_0_r[3 ] <= rom_data0[207:192]	;
			char_0_r[4 ] <= rom_data0[191:176]	;
			char_0_r[5 ] <= rom_data0[175:160]	;
			char_0_r[6 ] <= rom_data0[159:144]	;
			char_0_r[7 ] <= rom_data0[143:128]	;
			char_0_r[8 ] <= rom_data0[127:112]	;
			char_0_r[9 ] <= rom_data0[111:96]	;
			char_0_r[10] <= rom_data0[95:80]	;
			char_0_r[11] <= rom_data0[79:64]	;
			char_0_r[12] <= rom_data0[63:48]	;
			char_0_r[13] <= rom_data0[47:32]	;
			char_0_r[14] <= rom_data0[31:16]	;
			char_0_r[15] <= rom_data0[15:0]		;
		end
always@(posedge clk)
		begin
			char_1_r[0 ] <= rom_data1[255:240]	;
			char_1_r[1 ] <= rom_data1[239:224]	;
			char_1_r[2 ] <= rom_data1[223:208]	;
			char_1_r[3 ] <= rom_data1[207:192]	;
			char_1_r[4 ] <= rom_data1[191:176]	;
			char_1_r[5 ] <= rom_data1[175:160]	;
			char_1_r[6 ] <= rom_data1[159:144]	;
			char_1_r[7 ] <= rom_data1[143:128]	;
			char_1_r[8 ] <= rom_data1[127:112]	;
			char_1_r[9 ] <= rom_data1[111:96]	;
			char_1_r[10] <= rom_data1[95:80]	;
			char_1_r[11] <= rom_data1[79:64]	;
			char_1_r[12] <= rom_data1[63:48]	;
			char_1_r[13] <= rom_data1[47:32]	;
			char_1_r[14] <= rom_data1[31:16]	;
			char_1_r[15] <= rom_data1[15:0]		;
		end
always@(posedge clk)
		begin
			char_2_r[0 ] <= rom_data2[255:240]	;
			char_2_r[1 ] <= rom_data2[239:224]	;
			char_2_r[2 ] <= rom_data2[223:208]	;
			char_2_r[3 ] <= rom_data2[207:192]	;
			char_2_r[4 ] <= rom_data2[191:176]	;
			char_2_r[5 ] <= rom_data2[175:160]	;
			char_2_r[6 ] <= rom_data2[159:144]	;
			char_2_r[7 ] <= rom_data2[143:128]	;
			char_2_r[8 ] <= rom_data2[127:112]	;
			char_2_r[9 ] <= rom_data2[111:96]	;
			char_2_r[10] <= rom_data2[95:80]	;
			char_2_r[11] <= rom_data2[79:64]	;
			char_2_r[12] <= rom_data2[63:48]	;
			char_2_r[13] <= rom_data2[47:32]	;
			char_2_r[14] <= rom_data2[31:16]	;
			char_2_r[15] <= rom_data2[15:0]		;
        end
always@(posedge clk)
		begin
			char_3_r[0 ] <= rom_data3[255:240]	;
			char_3_r[1 ] <= rom_data3[239:224]	;
			char_3_r[2 ] <= rom_data3[223:208]	;
			char_3_r[3 ] <= rom_data3[207:192]	;
			char_3_r[4 ] <= rom_data3[191:176]	;
			char_3_r[5 ] <= rom_data3[175:160]	;
			char_3_r[6 ] <= rom_data3[159:144]	;
			char_3_r[7 ] <= rom_data3[143:128]	;
			char_3_r[8 ] <= rom_data3[127:112]	;
			char_3_r[9 ] <= rom_data3[111:96]	;
			char_3_r[10] <= rom_data3[95:80]	;
			char_3_r[11] <= rom_data3[79:64]	;
			char_3_r[12] <= rom_data3[63:48]	;
			char_3_r[13] <= rom_data3[47:32]	;
			char_3_r[14] <= rom_data3[31:16]	;
			char_3_r[15] <= rom_data3[15:0]		;
		end
always@(posedge clk)
		begin
			char_4_r[0 ] <= rom_data4[255:240]	;
			char_4_r[1 ] <= rom_data4[239:224]	;
			char_4_r[2 ] <= rom_data4[223:208]	;
			char_4_r[3 ] <= rom_data4[207:192]	;
			char_4_r[4 ] <= rom_data4[191:176]	;
			char_4_r[5 ] <= rom_data4[175:160]	;
			char_4_r[6 ] <= rom_data4[159:144]	;
			char_4_r[7 ] <= rom_data4[143:128]	;
			char_4_r[8 ] <= rom_data4[127:112]	;
			char_4_r[9 ] <= rom_data4[111:96]	;
			char_4_r[10] <= rom_data4[95:80]	;
			char_4_r[11] <= rom_data4[79:64]	;
			char_4_r[12] <= rom_data4[63:48]	;
			char_4_r[13] <= rom_data4[47:32]	;
			char_4_r[14] <= rom_data4[31:16]	;
			char_4_r[15] <= rom_data4[15:0]		;
		end
always@(posedge clk)
		begin
			char_5_r[0 ] <= rom_data5[255:240]	;
			char_5_r[1 ] <= rom_data5[239:224]	;
			char_5_r[2 ] <= rom_data5[223:208]	;
			char_5_r[3 ] <= rom_data5[207:192]	;
			char_5_r[4 ] <= rom_data5[191:176]	;
			char_5_r[5 ] <= rom_data5[175:160]	;
			char_5_r[6 ] <= rom_data5[159:144]	;
			char_5_r[7 ] <= rom_data5[143:128]	;
			char_5_r[8 ] <= rom_data5[127:112]	;
			char_5_r[9 ] <= rom_data5[111:96]	;
			char_5_r[10] <= rom_data5[95:80]	;
			char_5_r[11] <= rom_data5[79:64]	;
			char_5_r[12] <= rom_data5[63:48]	;
			char_5_r[13] <= rom_data5[47:32]	;
			char_5_r[14] <= rom_data5[31:16]	;
			char_5_r[15] <= rom_data5[15:0]		;
		end
always@(posedge clk)
		begin
			char_6_r[0 ] <= rom_data6[255:240]	;
			char_6_r[1 ] <= rom_data6[239:224]	;
			char_6_r[2 ] <= rom_data6[223:208]	;
			char_6_r[3 ] <= rom_data6[207:192]	;
			char_6_r[4 ] <= rom_data6[191:176]	;
			char_6_r[5 ] <= rom_data6[175:160]	;
			char_6_r[6 ] <= rom_data6[159:144]	;
			char_6_r[7 ] <= rom_data6[143:128]	;
			char_6_r[8 ] <= rom_data6[127:112]	;
			char_6_r[9 ] <= rom_data6[111:96]	;
			char_6_r[10] <= rom_data6[95:80]	;
			char_6_r[11] <= rom_data6[79:64]	;
			char_6_r[12] <= rom_data6[63:48]	;
			char_6_r[13] <= rom_data6[47:32]	;
			char_6_r[14] <= rom_data6[31:16]	;
			char_6_r[15] <= rom_data6[15:0]		;
		end
always@(posedge clk)
		begin
			char_7_r[0 ] <= rom_data7[255:240]	;
			char_7_r[1 ] <= rom_data7[239:224]	;
			char_7_r[2 ] <= rom_data7[223:208]	;
			char_7_r[3 ] <= rom_data7[207:192]	;
			char_7_r[4 ] <= rom_data7[191:176]	;
			char_7_r[5 ] <= rom_data7[175:160]	;
			char_7_r[6 ] <= rom_data7[159:144]	;
			char_7_r[7 ] <= rom_data7[143:128]	;
			char_7_r[8 ] <= rom_data7[127:112]	;
			char_7_r[9 ] <= rom_data7[111:96]	;
			char_7_r[10] <= rom_data7[95:80]	;
			char_7_r[11] <= rom_data7[79:64]	;
			char_7_r[12] <= rom_data7[63:48]	;
			char_7_r[13] <= rom_data7[47:32]	;
			char_7_r[14] <= rom_data7[31:16]	;
			char_7_r[15] <= rom_data7[15:0]		;
		end
always@(posedge clk)
		begin
			char_8_r[0 ] <= rom_data8[255:240]	;
			char_8_r[1 ] <= rom_data8[239:224]	;
			char_8_r[2 ] <= rom_data8[223:208]	;
			char_8_r[3 ] <= rom_data8[207:192]	;
			char_8_r[4 ] <= rom_data8[191:176]	;
			char_8_r[5 ] <= rom_data8[175:160]	;
			char_8_r[6 ] <= rom_data8[159:144]	;
			char_8_r[7 ] <= rom_data8[143:128]	;
			char_8_r[8 ] <= rom_data8[127:112]	;
			char_8_r[9 ] <= rom_data8[111:96]	;
			char_8_r[10] <= rom_data8[95:80]	;
			char_8_r[11] <= rom_data8[79:64]	;
			char_8_r[12] <= rom_data8[63:48]	;
			char_8_r[13] <= rom_data8[47:32]	;
			char_8_r[14] <= rom_data8[31:16]	;
			char_8_r[15] <= rom_data8[15:0]		;
		end
always@(posedge clk)
		begin
			char_9_r[0 ] <= rom_data9[255:240]	;
			char_9_r[1 ] <= rom_data9[239:224]	;
			char_9_r[2 ] <= rom_data9[223:208]	;
			char_9_r[3 ] <= rom_data9[207:192]	;
			char_9_r[4 ] <= rom_data9[191:176]	;
			char_9_r[5 ] <= rom_data9[175:160]	;
			char_9_r[6 ] <= rom_data9[159:144]	;
			char_9_r[7 ] <= rom_data9[143:128]	;
			char_9_r[8 ] <= rom_data9[127:112]	;
			char_9_r[9 ] <= rom_data9[111:96]	;
			char_9_r[10] <= rom_data9[95:80]	;
			char_9_r[11] <= rom_data9[79:64]	;
			char_9_r[12] <= rom_data9[63:48]	;
			char_9_r[13] <= rom_data9[47:32]	;
			char_9_r[14] <= rom_data9[31:16]	;
			char_9_r[15] <= rom_data9[15:0]		;
		end
endmodule
//    parameter bpos_x0=12'd180;
//    parameter bpos_y0=12'd360;
//   always@(*)
//         begin


//             if ( (Set_X>=bpos_x-12'd30) && (Set_X<=bpos_x+12'd30) )
//                begin
//                   if( (Set_Y>=bpos_y-12'd20) && (Set_Y<=bpos_y+12'd20) )
//                      RGB_Data<=24'h86edb0;
//                   else 
//                      begin
//                            if( Set_X >= pippos0_x1-12'd25 && Set_X <=pippos0_x1+12'd25 )
//                            begin
//                                  if( (Set_Y>=0 && Set_Y<=pippos0_y1)||( Set_Y>=pippos0_y2 && Set_Y<=12'd720 ) )
//                                  RGB_Data<= 24'h86c3ed;
//                                  else RGB_Data<=24'hffffff;
//                            end
//                            else RGB_Data<=24'hffffff;
//                      end
//                end
//             else if( Set_X >= pippos0_x1-12'd25 && Set_X <=pippos0_x1+12'd25 )
//               begin
//                   if( (Set_Y>=0 && Set_Y<=pippos0_y1)||( Set_Y>=pippos0_y2 && Set_Y<=12'd720 ) )
//                    RGB_Data<= 24'h86c3ed;
//                   else RGB_Data<=24'hffffff;
//               end
//             else
//                RGB_Data<=24'hffffff; 
//          end

//   always@(posedge clk)
//   begin
//     if(pos_y<=100) pos_y<=100;
//     else if(pos_y>=720) pos_y<=710;
//     else if(key1) pos_y<=pos_y+12'd2;
//     else if(key2) pos_y<=pos_y-12'd2;
//     else  pos_y<=pos_y; 
//   end

//    Picture_R_Rom R_ROM (
//      .clka(clk),    // input wire clka
//      .ena(1),      // input wire ena
//      .addra(Address),  // input wire [13 : 0] addra
//      .douta(R_Data)  // output wire [7 : 0] douta
//    );
//    Picture_G_Rom G_ROM (
//      .clka(clk),    // input wire clka
//      .ena(1),      // input wire ena
//      .addra(Address),  // input wire [13 : 0] addra
//      .douta(G_Data)  // output wire [7 : 0] douta
//    );
//    Picture_B_Rom B_ROM (
//      .clka(clk),    // input wire clka
//      .ena(1),      // input wire ena
//      .addra(Address),  // input wire [13 : 0] addra
//      .douta(B_Data)  // output wire [7 : 0] douta
//    );

// Number_Rom Number_Rom0(
//       .clka(clk),    // input wire clka
//       .ena(1),      // input wire ena
//       .addra(Address),  // input wire [13 : 0] addra
//       .douta(Num_Data)  // output wire [7 : 0] douta
// );
// else if(Set_X>=12'd1000&&Set_X<=12'd1015&&Set_Y>=12'd0&&Set_Y<=12'd15)
//     begin
//         Address=(Set_X-12'd999)*16+(Set_Y);
//         if(Num_Data) RGB_Data<=24'h0000ff;
//         else RGB_Data<=24'hffffff;
//     end

// else if(Set_X>=12'd1000&&Set_X<=12'd1015&&Set_Y>=12'd0&&Set_Y<=12'd15)
//     begin
//         if(char_5_r[Set_Y][12'd984-Set_X]) RGB_Data<=24'h20ffb2;
//         else RGB_Data<=24'hffbffa;
//     end
